module Demux(output [3:0]Y,input [1:0]A,input din);


    assign Y[0] = din & (~A[0]) & (~A[1]);
    assign Y[1] = din & (~A[1]) & A[0];
    assign Y[2] = din & A[1] & (~A[0]);
    assign Y[3] = din & A[1] & A[0];

endmodule